//Combining counter.sv and rom.sv:
//Counter module:
module counter#(
    parameter WIDTH = 8
)(

 // interface signals
 input logic [WIDTH-1:0] incr
 input logic clk, //input into counter block: clock
 input logic rst, //input into counter block: reset
 input logic en, //input into counter block: counter enable
 output logic [WIDTH-1:0] count //count output
);

always_ff @ (posedge clk)
    if (rst) count <= {WIDTH{1'b0}}; //so if rst is true (1) then count = 0
    else count<= count + {{WIDTH-1{1'b0}}, en}; //count increments by 1 as long as en is also true

endmodule

//ROM Module:
module rom # (
    parameter ADDRESS_WIDTH = 8, //Parameters are just the constants
              DATA_WIDTH = 8
)(
    //Assign input and output variables and their size:
    input logic clk,
    input logic [ADDRESS_WIDTH-1:0] addr, //address inputted into ROM is given by count of counter
    output logic [DATA_WIDTH-1:0] dout

);

//addr <= counter //so counter output is count which we assigned to addr

//Create 2D Array which is the ROM of size 2^8-1:0 (256 memory locations) and each memory location can hold 8-bit binary [7:0]
logic [DATA_WIDTH-1:0] rom_array [2**ADDRESS_WIDTH-1:0];

initial begin 
        $display("Loading rom.");
        $readmemh("sinerom.mem", rom_array); //sinerom.mem contains the data to store at the memory locations
        //sinerom.mem was generated by sinegen.py which goes through a cosine graph and inputs 256 of these values into a folder called sinerom.mem
        //these values are stored as hexadecimal
end;

always_ff @(posedge clk) 
    //So at positive clk edge, output the value at rom_array[addr]
    dout <= rom_array [addr]; 

endmodule

//Sinegen is 1 overall module that contains these 2 connected modules
module sinegen# (
  parameter WIDTH = 8
)

 // interface signals
 input logic [WIDTH-1:0] incr
 input logic clk, //input into singen block: clock
 input logic rst, //input into singen block: reset
 input logic en, //input into singen block: counter enable
 output logic [WIDTH-1:0] dout //singen output is the array output dout
);
//Similar to function calling in C++, input we send depends on what order inputs are initialized in modules and same for outputs

//Create variable which acts in the middle:
logic [WIDTH-1:0] addr //So this is what count from counter outputs to

counter firstCount (incr[7:0], clk, rst, en, addr[7:0]); //so instance of counter and output count is assigned to addr
rom lastRom (clk, addr[7:0], dout[7:0]); //so send inputs to ROM one of which is addr and assign output to dout[7:0];

endmodule

